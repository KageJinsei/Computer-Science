library verilog;
use verilog.vl_types.all;
entity turtle_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end turtle_vlg_check_tst;
