library verilog;
use verilog.vl_types.all;
entity turtle_vlg_vec_tst is
end turtle_vlg_vec_tst;
